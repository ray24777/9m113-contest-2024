module MatrixB (
    input   [127:0]   vsi_rdata,
    input   vsi_rdata_valid,
    output  [31:0]  
);
    
endmodule